module FPMUL_tb;
    initial begin
        $dumpfile("test.vcd");
        $dumpvars(0,test);  
    end
endmodule 