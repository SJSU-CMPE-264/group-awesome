`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// CMPE 140, CMPE Department, san Jose State University
// Authors: Donald Hung and Hoan Nguyen
//
// Create Date:    08:36:48 02/25/2010
// Design Name:
// Module Name:    mips_top
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
// MIPS Top-level Module (including the memories, clock,
// and the display module for prototyping)
module mips_top(
    input    clk, reset, pb,
    output    memwrite, wem, we1, we2, we3,
    output    [ 7:0]     LEDSEL,
    output     [ 7:0]    LEDOUT,
    input    [ 7:0]    switches,
    input   [7:0] gpi1,
    output    sinkBit
    
    );

    wire    [31:0]     pc, instr, dataadr, writedata, readdata, dispDat;
    wire    clksec, clk_db, faccel_done, FPM_done;
    reg     [ 15:0]    reg_hex;
    
    wire clk_5KHz;

    // Clock (1 second) to slow down the running of the instructions
    //clk_gen top_clk(.clk50MHz(clk), .reset(reset), .clksec(clksec));

    clk_gen top_clk(
        .clk100MHz(clk),
        .rst(reset),
        .clk_sec(clksec),
        .clk_5KHz(clk_5KHz)
        );
        
    debounce db (clk_5KHz, pb, clk_db);
      
    // Instantiate processor and memories    
    mips     mips       (clk_db, reset, pc, instr, memwrite, dataadr, writedata, readdata, switches[4:0], dispDat, (faccel_done | FPM_done));
    imem     imem       (pc[7:2], instr);
    //SoC
    SoC     soc ( 
                .addr(dataadr), .write_data(writedata), .gpi1(gpi1),
                .WE(memwrite), .reset(reset), .clk(clk_db), .data_out(readdata),
                .faccel_done(faccel_done), .FPM_done(FPM_done) 
                ); //faccel_done and FPM_done will be used for interrupt signal in full integration
    // decoder dec         (memwrite, dataadr, wem, we1, we2, we3, rdsel);
    // dmem    dmem        (clk_db, wem, dataadr, writedata, memdata);
    // faccel  fact        (clk_db, reset, we1, dataadr[3:2], writedata, fact_done_in, factdata);
    // gpio    gpio        (writedata, gpi1, 32'h0, dataadr[3:2], we2, clk_db, gpiodata, gpo1, gpo2);
    // FPWrapper FPWrapper (.clk(clk_db), .rst(reset), .A(dataadr[3:2]), .WE(we3), .InData(writedata), .done_sig(fp_done_in), .OutData(FPMdata));
    // register #(1) faccel_reg ( .clk(fact_done_in), .rst(dataadr[31:4] == fact_addr), .en(1'b1), .in(1'b1), .out(fact_done_out) );
    // register #(1) FP_reg ( .clk(fp_done_in), .rst(dataadr[31:4] == FP_addr), .en(1'b1), .in(1'b1), .out(fp_done_out) );
    // mux4 #(32) mux      (FPMdata, memdata, factdata, gpiodata, rdsel, readdata);
    
//=======================================================================================================================
//=======================================================================================================================

    wire [7:0] digit0;
    wire [7:0] digit1;
    wire [7:0] digit2;
    wire [7:0] digit3;
    wire [7:0] digit4;
    wire [7:0] digit5;
    wire [7:0] digit6;
    wire [7:0] digit7;
    
    bcd_to_7seg bcd0 (pc[15:12], digit0);
    bcd_to_7seg bcd1 (pc[11:8], digit1);
    bcd_to_7seg bcd2 (pc[7:4], digit2);
    bcd_to_7seg bcd3 (pc[3:0], digit3);
    
    bcd_to_7seg bcd4 (reg_hex[15:12], digit4);
    bcd_to_7seg bcd5 (reg_hex[11:8], digit5);
    bcd_to_7seg bcd6 (reg_hex[7:4], digit6);
    bcd_to_7seg bcd7 (reg_hex[3:0], digit7);
   
    LED_MUX disp_unit (
        clk_5KHz,
        reset,
        digit0,
        digit1,
        digit2,
        digit3,
        digit4,
        digit5,
        digit6,
        digit7,
        LEDOUT,
        LEDSEL        
        );
    
/*
    7:5 = 000 : Display LSW of register selected by DSW 4:0
    7:5 = 001 : Display MSW of register selected by DSW 4:0
    7:5 = 010 : Display LSW of instr
    7:5 = 011 : Display MSW of instr
    7:5 = 100 : DIsplay LSW of dataaddr
    7:5 = 101 : Display MSW of dataaddr
    7:5 = 110 : Display LSW of writedata
    7:5 = 111 : Display MSW of writedata
*/    
    
    always @ (posedge clk)
    begin
        case ({switches[7],switches[6], switches[5]})
            3'b000:    reg_hex = dispDat[15:0];
            3'b001:    reg_hex = dispDat[31:16];
            3'b010:    reg_hex = instr[15:0];
            3'b011:    reg_hex = instr[31:16];
            3'b100:    reg_hex = dataadr[15:0];
            3'b101:    reg_hex = dataadr[31:16];
            3'b110:    reg_hex = writedata[15:0];
            3'b111:    reg_hex = writedata[31:16];
            endcase
    end        

    //sink unused bit(s) to knock down the number of warning messages
    assign sinkBit = (pc > 0) ^ (instr > 0) ^ (dataadr > 0) ^ (writedata > 0) ^
                     (readdata > 0) ^ (dispDat > 0);
endmodule
